entity
library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;

  entity CTRL is
    port
      (
        
clk: in std logicvect
rst :in std_logic_vector
snd :in std_logic_vector
snd_led :out std_logic_vector

tx_data : out
tx_ready:
rx_data
rx_ready

baud_select
parity_select
